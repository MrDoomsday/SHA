`include "Ethalon/sha1.sv"